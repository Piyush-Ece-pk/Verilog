module moore_tb();
reg clk,rst,x;
wire z;

moore uut (
    .clk(clk),
    .rst(rst),
    .x(x),
    .z(z)
);

initial begin
    clk <= 1'b0;
    forever #5
    clk <= ~clk;
end

initial begin
    $dumpfile("dump.vcd");
    $dumpvars(0,moore_tb);
    rst <= 1'b0; #10;
    rst <= 1'b1;
    x <= 1'b1; #10;
    x <= 1'b1; #10;
    x <= 1'b1; #10;
    x <= 1'b0; #10;
    x <= 1'b1; #10;
    $finish;
end
endmodule

